// part1

module part1(
				clk
				);
	input logic clk;
endmodule